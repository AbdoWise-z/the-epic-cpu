Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

Entity Instruction_Mem is 

end Entity Instruction_Mem;


Architecture Instruction_Memarch of Instruction_Mem is
begin

end Architecture Instruction_Memarch;
