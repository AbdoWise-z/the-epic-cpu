entity StageDecode is
  port (
    clock
  ) ;
end StageDecode;