Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

Entity File_Register is 

end Entity File_Register;


Architecture File_Registerarch of File_Register is
begin

end Architecture File_Registerarch;
