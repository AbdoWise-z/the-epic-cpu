Library ieee;
use ieee.std_logic_1164.all;

Entity Forwarding_Unit is 

end Entity Forwarding_Unit;


Architecture Forwarding_Unitarch of Forwarding_Unit is
begin

end Architecture Forwarding_Unitarch;
