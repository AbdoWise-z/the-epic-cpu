Library ieee;
use ieee.std_logic_1164.all;

Entity ALU is 

end Entity ALU;


Architecture ALUarch of ALU is
begin

end Architecture ALUarch;