entity StageDecode is

end StageDecode;