Library ieee;
use ieee.std_logic_1164.all;

Entity Control_Unit is 

end Entity Control_Unit;


Architecture Control_Unitarch of Control_Unit is
begin
end Architecture Control_Unitarch;
