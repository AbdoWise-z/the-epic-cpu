Library ieee;
use ieee.std_logic_1164.all;

Entity Fetch is 

end Entity Fetch;


Architecture Fetcharch of Fetch is
begin

end Architecture Fetcharch;
